module hex_ssd (BIN, CLK, SSD);
	input [3:0] BIN;
	input CLK;
	output reg [0:6] SSD;
	
	always @(posedge CLK) begin
		case(BIN)
			0: SSD=7'b0000001;
			1: SSD=7'b1001111;
			2: SSD=7'b0010010;
			3: SSD=7'b0000110;
			4: SSD=7'b1001100;
			5: SSD=7'b0100100;
			6: SSD=7'b0100000;
			7: SSD=7'b0001111;
			8: SSD=7'b0000000;
			9: SSD=7'b0001100;
			10:SSD=7'b0001000;
			11:SSD=7'b1100000;
			12:SSD=7'b0110001;
			13:SSD=7'b1000010;
			14:SSD=7'b0110000;
			15:SSD=7'b0111000;
		endcase
	end
endmodule
